module not_gate


(input wire a,
output wire y);

assign y = ~a;

endmodule
